`define FD_BUS_Wid      32+1
`define DE_BUS_Wid      32+`alu_op_Wid+32+32+32+1+1+5+1
`define EM_BUS_Wid      32+32+1+5+1
`define MW_BUS_Wid      32+32+1+5
`define Branch_BUS_Wid  32+1
`define Wrf_BUS_Wid     32+1+5+32
`define ED_for_BUS_Wid  1+5+32
`define MD_for_BUS_Wid  5+32

`define alu_op_Wid      19

`define DCP0_BUS_Wid    
`define CP0D_BUS_Wid    
`define CP0E_BUS_Wid    
`define WCP0_BUS_Wid    